

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;
library gaisler;
use gaisler.misc.all;
library UNISIM;
use UNISIM.VComponents.all;


entity data_swapper is

 port(
 -- Clock and Reset -----------------
 HRDATA : out std_logic_vector (31 downto 0); -- AHB read-data
 dmao : in ahb_dma_out_type
 );
end;


architecture rtl of data_swapper is
begin
  HRDATA (7 downto 0) <= dmao.rdata(31 downto 24);
  HRDATA(15 downto 8) <= dmao.rdata(23 downto 16);
  HRDATA(23 downto 16) <= dmao.rdata(15 downto 8);
  HRDATA(31 downto 24) <= dmao.rdata(7 downto 0);
end;



